LIBRARY 	IEEE;
USE 		IEEE.STD_LOGIC_1164.ALL;
USE 		IEEE.NUMERIC_STD.all;

ENTITY ball_speed_rom IS
	PORT 
	(	
		diff_x		: IN	STD_LOGIC_VECTOR (2 DOWNTO 0);
		diff_y		: IN	STD_LOGIC_VECTOR (2 DOWNTO 0);
		speed_x		: OUT	STD_LOGIC_VECTOR (5 DOWNTO 0);
		speed_y		: OUT	STD_LOGIC_VECTOR (5 DOWNTO 0)
	);
END ball_speed_rom;

ARCHITECTURE behave OF ball_speed_rom IS

	TYPE rom_type IS ARRAY (0 TO 63) of UNSIGNED (5 DOWNTO 0);
	
	CONSTANT ROM_SPEED_X: rom_type :=
	(
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(20, 6),
		TO_UNSIGNED(15, 6),
		TO_UNSIGNED(12, 6),
		TO_UNSIGNED(10, 6),
		TO_UNSIGNED( 9, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(35, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(23, 6),
		TO_UNSIGNED(20, 6),
		TO_UNSIGNED(17, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(60, 6),
		TO_UNSIGNED(52, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(38, 6),
		TO_UNSIGNED(32, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(25, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(61, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(50, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(39, 6),
		TO_UNSIGNED(35, 6),
		TO_UNSIGNED(31, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED(58, 6),
		TO_UNSIGNED(54, 6),
		TO_UNSIGNED(49, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(40, 6),
		TO_UNSIGNED(37, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED(60, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(52, 6),
		TO_UNSIGNED(48, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(41, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED(61, 6),
		TO_UNSIGNED(58, 6),
		TO_UNSIGNED(55, 6),
		TO_UNSIGNED(51, 6),
		TO_UNSIGNED(48, 6),
		TO_UNSIGNED(45, 6)
	);

	CONSTANT ROM_SPEED_Y: rom_type :=
	(
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED(63, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(60, 6),
		TO_UNSIGNED(61, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED(62, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(52, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(58, 6),
		TO_UNSIGNED(60, 6),
		TO_UNSIGNED(61, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(20, 6),
		TO_UNSIGNED(35, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(50, 6),
		TO_UNSIGNED(54, 6),
		TO_UNSIGNED(56, 6),
		TO_UNSIGNED(58, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(15, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(38, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(49, 6),
		TO_UNSIGNED(52, 6),
		TO_UNSIGNED(55, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(12, 6),
		TO_UNSIGNED(23, 6),
		TO_UNSIGNED(32, 6),
		TO_UNSIGNED(39, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(48, 6),
		TO_UNSIGNED(51, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED(10, 6),
		TO_UNSIGNED(20, 6),
		TO_UNSIGNED(28, 6),
		TO_UNSIGNED(35, 6),
		TO_UNSIGNED(40, 6),
		TO_UNSIGNED(45, 6),
		TO_UNSIGNED(48, 6),
		TO_UNSIGNED( 0, 6),
		TO_UNSIGNED( 9, 6),
		TO_UNSIGNED(17, 6),
		TO_UNSIGNED(25, 6),
		TO_UNSIGNED(31, 6),
		TO_UNSIGNED(37, 6),
		TO_UNSIGNED(41, 6),
		TO_UNSIGNED(45, 6)
	);


BEGIN

	speed_x <= STD_LOGIC_VECTOR(ROM_SPEED_X(TO_INTEGER(UNSIGNED(diff_x & diff_y))));
	speed_y <= STD_LOGIC_VECTOR(ROM_SPEED_Y(TO_INTEGER(UNSIGNED(diff_x & diff_y))));

END behave;