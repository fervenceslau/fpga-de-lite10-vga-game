-- adc.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity adc is
	port (
		adc_pll_clock_clk        : in  std_logic                     := '0';             --  adc_pll_clock.clk
		adc_pll_locked_export    : in  std_logic                     := '0';             -- adc_pll_locked.export
		clock_clk                : in  std_logic                     := '0';             --          clock.clk
		command_valid            : in  std_logic                     := '0';             --        command.valid
		command_channel          : in  std_logic_vector(4 downto 0)  := (others => '0'); --               .channel
		command_startofpacket    : in  std_logic                     := '0';             --               .startofpacket
		command_endofpacket      : in  std_logic                     := '0';             --               .endofpacket
		command_ready            : out std_logic;                                        --               .ready
		command_2_valid          : in  std_logic                     := '0';             --      command_2.valid
		command_2_channel        : in  std_logic_vector(4 downto 0)  := (others => '0'); --               .channel
		command_2_startofpacket  : in  std_logic                     := '0';             --               .startofpacket
		command_2_endofpacket    : in  std_logic                     := '0';             --               .endofpacket
		command_2_ready          : out std_logic;                                        --               .ready
		reset_sink_reset_n       : in  std_logic                     := '0';             --     reset_sink.reset_n
		response_valid           : out std_logic;                                        --       response.valid
		response_channel         : out std_logic_vector(4 downto 0);                     --               .channel
		response_data            : out std_logic_vector(11 downto 0);                    --               .data
		response_startofpacket   : out std_logic;                                        --               .startofpacket
		response_endofpacket     : out std_logic;                                        --               .endofpacket
		response_2_valid         : out std_logic;                                        --     response_2.valid
		response_2_channel       : out std_logic_vector(4 downto 0);                     --               .channel
		response_2_data          : out std_logic_vector(11 downto 0);                    --               .data
		response_2_startofpacket : out std_logic;                                        --               .startofpacket
		response_2_endofpacket   : out std_logic                                         --               .endofpacket
	);
end entity adc;

architecture rtl of adc is
	component adc_modular_dual_adc_0 is
		port (
			clock_clk                : in  std_logic                     := 'X';             -- clk
			reset_sink_reset_n       : in  std_logic                     := 'X';             -- reset_n
			adc_pll_clock_clk        : in  std_logic                     := 'X';             -- clk
			adc_pll_locked_export    : in  std_logic                     := 'X';             -- export
			command_valid            : in  std_logic                     := 'X';             -- valid
			command_channel          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- channel
			command_startofpacket    : in  std_logic                     := 'X';             -- startofpacket
			command_endofpacket      : in  std_logic                     := 'X';             -- endofpacket
			command_ready            : out std_logic;                                        -- ready
			command_2_valid          : in  std_logic                     := 'X';             -- valid
			command_2_channel        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- channel
			command_2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			command_2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			command_2_ready          : out std_logic;                                        -- ready
			response_valid           : out std_logic;                                        -- valid
			response_channel         : out std_logic_vector(4 downto 0);                     -- channel
			response_data            : out std_logic_vector(11 downto 0);                    -- data
			response_startofpacket   : out std_logic;                                        -- startofpacket
			response_endofpacket     : out std_logic;                                        -- endofpacket
			response_2_valid         : out std_logic;                                        -- valid
			response_2_channel       : out std_logic_vector(4 downto 0);                     -- channel
			response_2_data          : out std_logic_vector(11 downto 0);                    -- data
			response_2_startofpacket : out std_logic;                                        -- startofpacket
			response_2_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component adc_modular_dual_adc_0;

begin

	modular_dual_adc_0 : component adc_modular_dual_adc_0
		port map (
			clock_clk                => clock_clk,                --          clock.clk
			reset_sink_reset_n       => reset_sink_reset_n,       --     reset_sink.reset_n
			adc_pll_clock_clk        => adc_pll_clock_clk,        --  adc_pll_clock.clk
			adc_pll_locked_export    => adc_pll_locked_export,    -- adc_pll_locked.export
			command_valid            => command_valid,            --        command.valid
			command_channel          => command_channel,          --               .channel
			command_startofpacket    => command_startofpacket,    --               .startofpacket
			command_endofpacket      => command_endofpacket,      --               .endofpacket
			command_ready            => command_ready,            --               .ready
			command_2_valid          => command_2_valid,          --      command_2.valid
			command_2_channel        => command_2_channel,        --               .channel
			command_2_startofpacket  => command_2_startofpacket,  --               .startofpacket
			command_2_endofpacket    => command_2_endofpacket,    --               .endofpacket
			command_2_ready          => command_2_ready,          --               .ready
			response_valid           => response_valid,           --       response.valid
			response_channel         => response_channel,         --               .channel
			response_data            => response_data,            --               .data
			response_startofpacket   => response_startofpacket,   --               .startofpacket
			response_endofpacket     => response_endofpacket,     --               .endofpacket
			response_2_valid         => response_2_valid,         --     response_2.valid
			response_2_channel       => response_2_channel,       --               .channel
			response_2_data          => response_2_data,          --               .data
			response_2_startofpacket => response_2_startofpacket, --               .startofpacket
			response_2_endofpacket   => response_2_endofpacket    --               .endofpacket
		);

end architecture rtl; -- of adc
